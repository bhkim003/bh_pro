module{

}
endmodule
